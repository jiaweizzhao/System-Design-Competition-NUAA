`timescale 1ns / 1ps
//*************************************************************************
//   > �ļ���: decode.v
//   > ����  :�弶��ˮCPU������ģ��
//   > ����  : LOONGSON
//   > ����  : 2016-04-14
//*************************************************************************
module decode(                      // ���뼶
    input              ID_valid,    // ���뼶��Ч�ź�
    input      [ 63:0] IF_ID_bus_r, // IF->ID����
    input      [ 31:0] rs_value,    // ��һԴ������ֵ
    input      [ 31:0] rt_value,    // �ڶ�Դ������ֵ
    output     [  4:0] rs,          // ��һԴ��������ַ 
    output     [  4:0] rt,          // �ڶ�Դ��������ַ
    output     [ 32:0] jbr_bus,     // ��ת����
//  output             inst_jbr,    // ָ��Ϊ��ת��ָ֧��,�弶��ˮ����Ҫ
    output             ID_over,     // IDģ��ִ�����
    output     [202:0] ID_EXE_bus,  // ID->EXE����
    
    //5����ˮ����
    input              IF_over,     //���ڷ�ָ֧���Ҫ���ź�
    input      [  4:0] EXE_wdest,   // EXE��Ҫд�ؼĴ����ѵ�Ŀ���ַ��
    input      [  4:0] MEM_wdest,   // MEM��Ҫд�ؼĴ����ѵ�Ŀ���ַ��
    input      [  4:0] WB_wdest,    // WB��Ҫд�ؼĴ����ѵ�Ŀ���ַ��
    

    input             cal_r_E,
    input             cal_i_E,
    input             lui_E,
    input             mf_E,
    input             load_E,
    input             mf_M,
    input             load_M,
    input             Q,
    //չʾPC
    output     [ 31:0] ID_pc
);
//-----{IF->ID����}begin
    wire [31:0] pc;
    wire [31:0] inst;
    assign {pc, inst} = IF_ID_bus_r;  // IF->ID���ߴ�PC��ָ��
//-----{IF->ID����}end

//-----{ָ������}begin
    wire [5:0] op;       
    wire [4:0] rd;       
    wire [4:0] sa;      
    wire [5:0] funct;    
    wire [15:0] imm;     
    wire [15:0] offset;  
    wire [25:0] target;  
    wire [2:0] cp0r_sel;

    assign op     = inst[31:26];  // ������
    assign rs     = inst[25:21];  // Դ������1
    assign rt     = inst[20:16];  // Դ������2
    assign rd     = inst[15:11];  // Ŀ�������
    assign sa     = inst[10:6];   // �����򣬿��ܴ��ƫ����
    assign funct  = inst[5:0];    // ������
    assign imm    = inst[15:0];   // ������
    assign offset = inst[15:0];   // ��ַƫ����
    assign target = inst[25:0];   // Ŀ���ַ
    assign cp0r_sel= inst[2:0];   // cp0�Ĵ�����select��

    // ʵ��ָ���б�
    wire inst_ADDU, inst_SUBU , inst_SLT , inst_AND;
    wire inst_ADD , inst_SUB  , inst_ADDI, inst_DIV;
    wire inst_NOR , inst_OR   , inst_XOR , inst_SLL;
    wire inst_SRL , inst_ADDIU, inst_BEQ , inst_BNE;
    wire inst_LW  , inst_SW   , inst_LUI , inst_J;
    wire inst_SLTU, inst_JALR , inst_JR  , inst_SLLV;
    wire inst_SRA , inst_SRAV , inst_SRLV, inst_SLTIU;
    wire inst_SLTI, inst_BGEZ , inst_BGTZ, inst_BLEZ;
    wire inst_BLTZ, inst_LB   , inst_LBU , inst_SB;
    wire inst_ANDI, inst_ORI  , inst_XORI, inst_JAL;
    wire inst_MULT, inst_MFLO , inst_MFHI, inst_MTLO;
    wire inst_MTHI, inst_MFC0 , inst_MTC0;
    wire inst_MULTU, inst_DIVU;
    wire inst_LH, inst_LHU, inst_SH;
    wire inst_ERET, inst_SYSCALL, inst_BREAK;
    wire inst_BLTZAL, inst_BGEZAL;


    wire op_zero;  // ������ȫ0
    wire sa_zero;  // sa��ȫ0
    assign op_zero = ~(|op);
    assign sa_zero = ~(|sa);
    assign inst_ADDU  = op_zero & sa_zero    & (funct == 6'b100001);//�޷��żӷ�
    assign inst_SUBU  = op_zero & sa_zero    & (funct == 6'b100011);//�޷��ż���
    assign inst_ADD   = op_zero & sa_zero    & (funct == 6'b100000);//�з��żӷ�
    assign inst_SUB   = op_zero & sa_zero    & (funct == 6'b100010);//�з��ż���
    assign inst_SLT   = op_zero & sa_zero    & (funct == 6'b101010);//С������λ
    assign inst_SLTU  = op_zero & sa_zero    & (funct == 6'b101011);//�޷���С����
    assign inst_JALR  = op_zero & (rt==5'd0) & (rd==5'd31)
                      & sa_zero & (funct == 6'b001001);         //��ת�Ĵ���������
    assign inst_JR    = op_zero & (rt==5'd0) & (rd==5'd0 )
                      & sa_zero & (funct == 6'b001000);             //��ת�Ĵ���
    assign inst_AND   = op_zero & sa_zero    & (funct == 6'b100100);//������
    assign inst_NOR   = op_zero & sa_zero    & (funct == 6'b100111);//�������
    assign inst_OR    = op_zero & sa_zero    & (funct == 6'b100101);//������
    assign inst_XOR   = op_zero & sa_zero    & (funct == 6'b100110);//�������
    assign inst_SLL   = op_zero & (rs==5'd0) & (funct == 6'b000000);//�߼�����
    assign inst_SLLV  = op_zero & sa_zero    & (funct == 6'b000100);//�����߼�����
    assign inst_SRA   = op_zero & (rs==5'd0) & (funct == 6'b000011);//��������
    assign inst_SRAV  = op_zero & sa_zero    & (funct == 6'b000111);//������������
    assign inst_SRL   = op_zero & (rs==5'd0) & (funct == 6'b000010);//�߼�����
    assign inst_SRLV  = op_zero & sa_zero    & (funct == 6'b000110);//�����߼�����
    assign inst_MULT  = op_zero & (rd==5'd0)
                      & sa_zero & (funct == 6'b011000);             //�˷�
    assign inst_MULTU  = op_zero & (rd==5'd0)
                      & sa_zero & (funct == 6'b011001);             //�޷������˷�
    assign inst_DIV   = op_zero & (rd==5'd0)
                      & sa_zero & (funct == 6'b011010);             //����
    assign inst_DIVU  = op_zero & (rd==5'd0)
                      & sa_zero & (funct == 6'b011011);             //�޷��ų���               
    assign inst_MFLO  = op_zero & (rs==5'd0) & (rt==5'd0)
                      & sa_zero & (funct == 6'b010010);             //��LO��ȡ
    assign inst_MFHI  = op_zero & (rs==5'd0) & (rt==5'd0)
                      & sa_zero & (funct == 6'b010000);             //��HI��ȡ
    assign inst_MTLO  = op_zero & (rt==5'd0) & (rd==5'd0)
                      & sa_zero & (funct == 6'b010011);             //��LOд����
    assign inst_MTHI  = op_zero & (rt==5'd0) & (rd==5'd0)
                      & sa_zero & (funct == 6'b010001);             //��HIд����
    assign inst_ADDIU = (op == 6'b001001);             //�������޷��żӷ�
    assign inst_ADDI  = (op == 6'b001000);			   //�������ӷ�
    assign inst_SLTI  = (op == 6'b001010);             //С������������λ
    assign inst_SLTIU = (op == 6'b001011);             //С������������λ���޷��ţ�
    assign inst_BEQ   = (op == 6'b000100);             //�ж������ת
    assign inst_BGEZ  = (op == 6'b000001) & (rt==5'd1);//���ڵ���0��ת
    assign inst_BGTZ  = (op == 6'b000111) & (rt==5'd0);//����0��ת
    assign inst_BLEZ  = (op == 6'b000110) & (rt==5'd0);//С�ڵ���0��ת
    assign inst_BLTZ  = (op == 6'b000001) & (rt==5'd0);//С��0��ת
    assign inst_BNE   = (op == 6'b000101);             //�жϲ�����ת
    assign inst_LW    = (op == 6'b100011);             //���ڴ�װ����
    assign inst_SW    = (op == 6'b101011);             //���ڴ�洢��
    assign inst_LB    = (op == 6'b100000);             //load�ֽڣ�������չ��
    assign inst_LBU   = (op == 6'b100100);             //load�ֽڣ��޷�����չ��
    assign inst_SB    = (op == 6'b101000);             //���ڴ�洢�ֽ�
    assign inst_LH    = (op == 6'b100001);             //���ڴ�װ�ذ��֣�������չ��
    assign inst_LHU   = (op == 6'b100101);             //���ڴ�װ�ذ��֣��޷�����չ��
    assign inst_SH    = (op == 6'b101001);             //���ڴ�洢��
    assign inst_ANDI  = (op == 6'b001100);             //��������
    assign inst_LUI   = (op == 6'b001111) & (rs==5'd0);//������װ�ظ߰��ֽ�
    assign inst_ORI   = (op == 6'b001101);             //��������
    assign inst_XORI  = (op == 6'b001110);             //���������
    assign inst_J     = (op == 6'b000010);             //��ת
    assign inst_JAL   = (op == 6'b000011);             //��ת������
    assign inst_MFC0    = (op == 6'b010000) & (rs==5'd0) 
                        & sa_zero & (funct[5:3] == 3'b000); // ��cp0�Ĵ���װ��
    assign inst_MTC0    = (op == 6'b010000) & (rs==5'd4)
                        & sa_zero & (funct[5:3] == 3'b000); // ��cp0�Ĵ����洢
    assign inst_SYSCALL = (op == 6'b000000) & (funct == 6'b001100); // ϵͳ����
    assign inst_ERET    = (op == 6'b010000) & (rs==5'd16) & (rt==5'd0)
                        & (rd==5'd0) & sa_zero & (funct == 6'b011000);//�쳣����

    assign inst_BREAK  = (op == 6'b000000) & (funct == 6'b001101); //�����ϵ�����

    assign inst_BLTZAL = (op == 6'b000001)& (rt==5'b10000);//С������ת����31�żĴ�������
    assign inst_BGEZAL = (op == 6'b000001)& (rt==5'b10001);//���ڵ�������ת����31�żĴ�������
            
            //ȱ��break bltzal bgezal�Ķ���
    
    //��ת��ָ֧��
    wire inst_jr;    //�Ĵ�����תָ��
    wire inst_j_link;//������תָ��
    wire inst_jbr;   //���з�֧��תָ��
    assign inst_jr     = inst_JALR | inst_JR;
    assign inst_j_link = inst_JAL | inst_JALR |inst_BLTZAL | inst_BGEZAL;
    assign inst_jbr = inst_J    | inst_JAL  | inst_jr
                    | inst_BEQ  | inst_BNE  | inst_BGEZ
                    | inst_BGTZ | inst_BLEZ | inst_BLTZ
                    | inst_BLTZAL | inst_BGEZAL;
        
    //load store
    wire inst_load;
    wire inst_store;
    assign inst_load  = inst_LW | inst_LB | inst_LBU | inst_LH | inst_LHU;  // loadָ��
    assign inst_store = inst_SW | inst_SB | inst_SH;                        // storeָ��
    
    //alu��������
    wire inst_add, inst_sub, inst_slt,inst_sltu;
    wire inst_and, inst_nor, inst_or, inst_xor;
    wire inst_sll, inst_srl, inst_sra,inst_lui;
    wire inst_overflow;

    assign inst_add = inst_ADDU | inst_ADDIU | inst_load
                    | inst_store | inst_j_link |inst_ADD
                    | inst_ADDI; 			              // ���ӷ�
    assign inst_sub = inst_SUBU | inst_SUB;                // ����
    assign inst_slt = inst_SLT | inst_SLTI;                // �з���С����λ
    assign inst_sltu= inst_SLTIU | inst_SLTU;              // �޷���С����λ
    assign inst_and = inst_AND | inst_ANDI;                // �߼���
    assign inst_nor = inst_NOR;                            // �߼����
    assign inst_or  = inst_OR  | inst_ORI;                 // �߼���
    assign inst_xor = inst_XOR | inst_XORI;                // �߼����
    assign inst_sll = inst_SLL | inst_SLLV;                // �߼�����
    assign inst_srl = inst_SRL | inst_SRLV;                // �߼�����
    assign inst_sra = inst_SRA | inst_SRAV;                // ��������
    assign inst_lui = inst_LUI;                            // ������װ�ظ�λ
    assign inst_overflow = inst_ADDI | inst_ADD |inst_SUB; // �з������
    
    //ʹ��sa����Ϊƫ��������λָ��
    wire inst_shf_sa;
    assign inst_shf_sa =  inst_SLL | inst_SRL | inst_SRA;
    
    //������������չ��ʽ����
    wire inst_imm_zero; //������0��չ
    wire inst_imm_sign; //������������չ
    assign inst_imm_zero = inst_ANDI  | inst_LUI  | inst_ORI | inst_XORI;
    assign inst_imm_sign = inst_ADDIU |  inst_SLTI | inst_SLTIU
                         | inst_load | inst_store | inst_ADDI;
    
    //����Ŀ�ļĴ����ŷ���
    wire inst_wdest_rt;  // �Ĵ�����д���ַΪrt��ָ��
    wire inst_wdest_31;  // �Ĵ�����д���ַΪ31��ָ��  
    wire inst_wdest_rd;  // �Ĵ�����д���ַΪrd��ָ��
    assign inst_wdest_rt = inst_imm_zero | inst_ADDIU | inst_SLTI | inst_ADDI
                         | inst_SLTIU | inst_load | inst_MFC0;
    assign inst_wdest_31 = inst_JAL |inst_BLTZAL | inst_BGEZAL;
    assign inst_wdest_rd = inst_ADDU | inst_SUBU | inst_SLT  | inst_SLTU
                         | inst_JALR | inst_AND  | inst_NOR  | inst_OR 
                            | inst_XOR  | inst_SLL  | inst_SLLV | inst_SRA 
                         | inst_SRAV | inst_SRL  | inst_SRLV
                         | inst_MFHI | inst_MFLO | inst_ADD | inst_SUB;
                         
    //����Դ�Ĵ����ŷ���
    wire inst_no_rs;  //ָ��rs���0���Ҳ��ǴӼĴ����Ѷ�rs������
    wire inst_no_rt;  //ָ��rt���0���Ҳ��ǴӼĴ����Ѷ�rt������
    assign inst_no_rs = inst_MTC0 | inst_SYSCALL | inst_ERET | inst_BREAK;
    assign inst_no_rt = inst_ADDIU | inst_SLTI | inst_SLTIU
                      | inst_BGEZ  | inst_load | inst_imm_zero
                      | inst_J     | inst_JAL  | inst_MFC0
                      | inst_SYSCALL | inst_ADDI |inst_BLTZAL | inst_BGEZAL | inst_BREAK;
//-----{ָ������}end

//-----{��ָ֧��ִ��}begin
   //bd_pc,��֧��תָ���������Ϊ�ӳٲ�ָ���PCֵ������ǰ��ָ֧���PC+4
    wire [31:0] bd_pc;   //�ӳٲ�ָ��PCֵ
    assign bd_pc = pc + 3'b100;
    
    //��������ת
    wire        j_taken;
    wire [31:0] j_target;
    assign j_taken = inst_J | inst_JAL | inst_jr;
    //�Ĵ�����ת��ַΪrs_value,������תΪ{bd_pc[31:28],target,2'b00}
    assign j_target = inst_jr ? rs_value : {bd_pc[31:28],target,2'b00};

    //branchָ��
    wire rs_equql_rt;
    wire rs_ez;
    wire rs_ltz;
    assign rs_equql_rt = (rs_value == rt_value);  // GPR[rs]==GPR[rt]
    assign rs_ez       = ~(|rs_value);            // rs�Ĵ���ֵΪ0
    assign rs_ltz      = rs_value[31];            // rs�Ĵ���ֵС��0
    wire br_taken;
    wire [31:0] br_target;
    assign br_taken = inst_BEQ  & rs_equql_rt       // �����ת
                    | inst_BNE  & ~rs_equql_rt      // ������ת
                    | (inst_BGEZ | inst_BGEZAL) & ~rs_ltz           // ���ڵ���0��ת
                    | inst_BGTZ & ~rs_ltz & ~rs_ez  // ����0��ת
                    | inst_BLEZ & (rs_ltz | rs_ez)  // С�ڵ���0��ת
                    | (inst_BLTZ | inst_BLTZAL) & rs_ltz;           // С��0��ת
    // ��֧��תĿ���ַ��PC=PC+offset<<2
    assign br_target[31:2] = bd_pc[31:2] + {{14{offset[15]}}, offset};  
    assign br_target[1:0]  = bd_pc[1:0];
    
    //jump and branchָ��
    wire jbr_taken;
    wire [31:0] jbr_target;
    assign jbr_taken = (j_taken | br_taken) & ID_over; 
    assign jbr_target = j_taken ? j_target : br_target;
    
    //ID��IF����ת����
    assign jbr_bus = {jbr_taken, jbr_target};
//-----{��ָ֧��ִ��}end

//-----{IDִ�����}begin
    //��������ˮ�ģ������������
    //wire rs_wait;
    //wire rt_wait;
    /*assign rs_wait = ~inst_no_rs & (rs!=5'd0)
                   & ( (rs==EXE_wdest) | (rs==MEM_wdest) | (rs==WB_wdest) );
    assign rt_wait = ~inst_no_rt & (rt!=5'd0)
                   & ( (rt==EXE_wdest) | (rt==MEM_wdest) | (rt==WB_wdest) );*/
    
    //���ڷ�֧��תָ�ֻ����IFִ����ɺ󣬲ſ�����ID��ɣ�
    //����ID��������ˣ���IF����ȡָ���next_pc�������浽PC��ȥ��
    //��ô��IF��ɣ�next_pc�����浽PC��ȥʱ��jbr_bus�ϵ������ѱ����Ч��
    //���·�֧��תʧ��
    //(~inst_jbr | IF_over)����(~inst_jbr | (inst_jbr & IF_over))
    assign ID_over = ID_valid & stall & (~inst_jbr | IF_over);
//-----{IDִ�����}end

//-----{ID->EXE����}begin
    //���������ʵ�Ǽ���ʽ��ֲ�ʽ��ϵ�˼�룬��Ȼ�źŶ���ID�׶����ɣ��������ɵ�ÿ���ź�ֻ��һ���׶�ʹ�ã����źŰ��׶����ֿ�����Ȼ��ÿ���׶��л����źŵ�����
    //EXE��Ҫ�õ�����Ϣ
    wire multiply;         //�˷�MULT
    wire divide;           //����DIV
    wire sign_exe;         //�˳������޷������ж�
    wire mthi;             //MTHI
    wire mtlo;             //MTLO
    assign multiply = inst_MULT | inst_MULTU;
    assign divide = inst_DIV | inst_DIVU;
    assign sign_exe = inst_MULT | inst_DIV;
    assign mthi     = inst_MTHI ;
    assign mtlo     = inst_MTLO;

    //ALU����Դ�������Ϳ����ź�
    wire [12:0] alu_control;
    wire [31:0] alu_operand1;
    wire [31:0] alu_operand2;
    
    //��ν������ת�ǽ���ת���ص�PCֵ��ŵ�31�żĴ�����
    //����ˮCPU������ӳٲۣ���������ת��Ҫ����PC+8����ŵ�31�żĴ�����
    assign alu_operand1 = inst_j_link ? pc : 
                          inst_shf_sa ? {27'd0,sa} : rs_value;
    assign alu_operand2 = inst_j_link ? 32'd8 :  
                          inst_imm_zero ? {16'd0, imm} :
                          inst_imm_sign ?  {{16{imm[15]}}, imm} : rt_value;
    assign alu_control = {inst_overflow,    // ALU�����룬���ȱ���
                          inst_add,        
                          inst_sub,
                          inst_slt,
                          inst_sltu,
                          inst_and,
                          inst_nor,
                          inst_or, 
                          inst_xor,
                          inst_sll,
                          inst_srl,
                          inst_sra,
                          inst_lui
                          };

    //�ô���Ҫ�õ���load/store��Ϣ
    wire       lb_sign;  //loadһ�ֽ�Ϊ�з���load
    wire       lh_sign;  //load����Ϊ�з���load
    wire [1:0] ls_word;  //load/storeΪ�ֽڻ����ֻ��ǰ���,00:byte;10:word;half:01
    wire [5:0] mem_control;  //MEM��Ҫʹ�õĿ����ź�
    wire [31:0] store_data;  //store�����Ĵ������
    assign lb_sign = inst_LB ;
    assign lh_sign = inst_LH ;
    assign ls_word = {inst_LW | inst_SW, inst_LH | inst_SH};
    assign mem_control = {inst_load,
                          inst_store,
                          ls_word,
                          lb_sign,
                          lh_sign};
                          
    //д����Ҫ�õ�����Ϣ
    wire mfhi;
    wire mflo;
    wire mtc0;
    wire mfc0;
    wire [7 :0] cp0r_addr;
    wire       syscall;   //syscall��eret��д�ؼ�������Ĳ��� 
    wire       eret;
    wire       rf_wen;    //д�صļĴ���дʹ��
    wire [4:0] rf_wdest;  //д�ص�Ŀ�ļĴ���
    assign syscall  = inst_SYSCALL;
    assign break    = inst_BREAK;//����һ������break�Ŀ����ź�
    assign eret     = inst_ERET;
    assign mfhi     = inst_MFHI;
    assign mflo     = inst_MFLO;
    assign mtc0     = inst_MTC0;
    assign mfc0     = inst_MFC0;
    assign cp0r_addr= {rd,cp0r_sel};
    assign rf_wen   = inst_wdest_rt | inst_wdest_31 | inst_wdest_rd;
    assign rf_wdest = inst_wdest_rt ? rt :     //�ڲ�д�Ĵ�����ʱ����Ϊ0
                      inst_wdest_31 ? 5'd31 :  //�Ա���׼ȷ�ж��������
                      inst_wdest_rd ? rd : 5'd0;
    assign store_data = rt_value;
    assign ID_EXE_bus = {
                         outsa,
                         inst_j_link,
                         rs,rt,rd,
                         cal_r_D,cal_i_D,store_D,load_D,jump_D,mt_D,CMPOp, ID_b_type,ID_b_zero,
                         mf_D,lui_D,
                         multiply,divide,sign_exe,mthi,mtlo,   //EXE���õ���Ϣ,����
                         alu_control,alu_operand1,alu_operand2,//EXE���õ���Ϣ
                         mem_control,store_data,               //MEM���õ��ź�
                         mfhi,mflo,                            //WB���õ��ź�,����
                         mtc0,mfc0,cp0r_addr,syscall,break,eret,     //WB���õ��ź�,����
                         rf_wen, rf_wdest,                     //WB���õ��ź�
                         pc                                   //PCֵ
                        };    

//-----{ID->EXE����}end

//-----{չʾIDģ���PCֵ}begin
    assign ID_pc = pc;
//-----{չʾIDģ���PCֵ}end

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//stallģ��
wire stall;
wire stall_cal_r;
wire stall_cal_i;
wire stall_beq;
wire stall_jump;
wire stall_load;
wire stall_store;
wire stall_mt;

wire cal_r_D;
wire cal_i_D;
wire store_D;
wire load_D;
wire jump_D;
wire mt_D;
wire beq_D;
wire mf_D;
wire lui_D;

wire ID_b_type;
wire ID_b_zero;
wire [4:0] outsa;
wire sl;

assign sl = inst_sll | inst_srl | inst_sra ;
assign jump_D = inst_jr;
assign cal_r_D = inst_ADD | inst_ADDU | inst_SUB |inst_SUBU |inst_SLTU | inst_SLT | inst_DIV |inst_DIVU | inst_MULT | inst_MULTU | inst_AND |inst_NOR |inst_OR | inst_XOR | inst_SLLV |inst_SLL |inst_SRAV |inst_SRA | inst_SRLV |inst_SRL;
assign cal_i_D = inst_ADDI | inst_ADDIU | inst_SLTIU | inst_SLTI | inst_ANDI |inst_ORI | inst_XORI;
assign beq_D = inst_BEQ | inst_BNE |inst_BGEZ |inst_BGTZ |inst_BLEZ |inst_BLTZ |inst_BGEZAL |inst_BLTZAL;
assign load_D = inst_LB | inst_LBU | inst_LH |inst_LHU |inst_LW;
assign store_D = inst_SB |inst_SH |inst_SW;
assign mt_D = inst_MTHI |inst_MTLO ;
assign lui_D = inst_LUI;
assign mf_D = inst_MFLO | inst_MFHI;
assign ID_b_type = inst_BEQ | inst_BNE;
assign ID_b_zero = inst_BGEZ | inst_BGTZ |inst_BLEZ |inst_BLTZ |inst_BGEZAL |inst_BLTZAL;

assign stall_beq = beq_D & ( (cal_r_E & ((rs == EXE_wdest) | (rt == EXE_wdest))) | 
                             (cal_i_E & ((rs == EXE_wdest) | (rt == EXE_wdest))) | 
                             (lui_E   & ((rs == EXE_wdest) | (rt == EXE_wdest))) |
                             (mf_E    & ((rs == EXE_wdest) | (rt == EXE_wdest))) | 
                             (load_E  & ((rs == EXE_wdest) | (rt == EXE_wdest))) |
                             (mf_M    & ((rs == MEM_wdest) | (rt == MEM_wdest))) |
                             (load_M  & ((rs == MEM_wdest) | (rt == MEM_wdest)))
                           );

assign stall_cal_r  = cal_r_D & (
                                  (mf_E    & ((rs == EXE_wdest) | (rt == EXE_wdest))) |
                                  (load_E  & ((rs == EXE_wdest) | (rt == EXE_wdest))) 
                                ); 
assign stall_cal_i  = cal_i_D & (
                                  (mf_E    & (rs == EXE_wdest)) |
                                  (load_E  & (rs == EXE_wdest)) 
                                );
assign stall_load   = load_D  & (
                                  (mf_E    & (rs == EXE_wdest)) |
                                  (load_E  & (rs == EXE_wdest))    
                                );
assign stall_store  = store_D & (
                                  (mf_E    & (rs == EXE_wdest)) |
                                  (load_E  & (rs == EXE_wdest))    
                                );
assign stall_jump   = jump_D  & (
                                    (cal_r_E & (rs == EXE_wdest)) | 
                                    (cal_i_E & (rs == EXE_wdest)) | 
                                    (lui_E   & (rs == EXE_wdest)) |
                                    (mf_E    & (rs == EXE_wdest)) | 
                                    (load_E  & (rs == EXE_wdest)) |
                                    (mf_M    & (rs == MEM_wdest)) |
                                    (load_M  & (rs == MEM_wdest))
                                );
assign  stall_mt    = mt_D    & (
                                    (cal_r_E & (rs == EXE_wdest)) | 
                                    (cal_i_E & (rs == EXE_wdest)) | 
                                    (lui_E   & (rs == EXE_wdest)) |
                                    (mf_E    & (rs == EXE_wdest)) | 
                                    (load_E  & (rs == EXE_wdest)) |
                                    (mf_M    & (rs == MEM_wdest)) |
                                    (load_M  & (rs == MEM_wdest))
                                );
assign stall =  stall_cal_r | stall_cal_i | stall_beq | stall_jump | stall_load | stall_store | stall_mt;

assign outsa =  (sl) ? sa : 5'b0;
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

assign CMPOp =  inst_BEQ  ? 3'b000 :
                inst_BNE  ? 3'b001 :
                inst_BLEZ ? 3'b010 :
                inst_BGTZ ? 3'b011 :
                inst_BLTZ ? 3'b100 :
                inst_BGEZ ? 3'b101 :
                inst_BLTZAL? 3'b110:
                inst_BGEZAL? 3'b111;
wire PCSel;
wire Flush;

assign PCSel = ( inst_jr  )                                 ? 2 :
               ( inst_J    ||  inst_JAL ||  (beq_D && Q ))  ? 1 : 
                                                              0 ;
assign Flush = (PCSel == 1)||(PCSel == 2);




endmodule
